/*
This is a useless file.
*/