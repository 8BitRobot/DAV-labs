module miniALU(
	/* TODO: Ports go here (refer to lab spec) */
);
	// The following block will contain the logic of your combinational circuit
	always_comb begin
		/* TODO: Depending on the value of your select bit, output the result of a different operation.
		 * Refer to the lab spec for details. 
		 */
	end
endmodule