module miniALU(
	/* Ports go here */
);

	// The following block will contain the logic of your combinational circuit
	always_comb begin
		/* How can you set result to a different value depending on the value of
		   your select line? */
	end
endmodule