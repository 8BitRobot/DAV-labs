module fft (
	
);



endmodule