module alarmClock_top (
input PSS_button, input reset_button, input clk, input [5:0] time_switches, input speed_switch, 
output logic [7:0] display [5:0]
);


endmodule