
//TODO: Finish nunchuck_translator as described in the lab spec!