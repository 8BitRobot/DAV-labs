module nunchuck_test(clk, rst, sda, scl);
	
	//TODO: Modify this file to do something meaningful with the nunchuck!
	
	
endmodule