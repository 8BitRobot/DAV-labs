`timescale 1ns/1ns

module twiddle_module 
(
	input clk,
	input [3:0] stage, 
	input [9:0] address_a,
	output reg [47:00] twiddle
);

	wire [9:0] select_raw;
	wire [8:0] select;
	
	assign select_raw = address_a << (4'b1001 - stage);
	assign select = select_raw[8:0];
	
	manual_twiddle_rom twiddle_rom(
		.address(select),
		.clock(clk),
		.q(twiddle)
	);
	
endmodule 

module manual_twiddle_rom (
	input [8:0] address,
	input clock,
	output reg [47:00] q
);


	always @(posedge clock) begin
		case (address)
		
			  0: q = 48'h7FFFFF000000;
			  1: q = 48'h7FFF6200C910;
			  2: q = 48'h7FFD8801921D;
			  3: q = 48'h7FFA73025B27;
			  4: q = 48'h7FF62203242B;
			  5: q = 48'h7FF09403ED27;
			  6: q = 48'h7FE9CC04B619;
			  7: q = 48'h7FE1C7057F00;
			  8: q = 48'h7FD8880647D9;
			  9: q = 48'h7FCE0C0710A3;
			 10: q = 48'h7FC25607D95C;
			 11: q = 48'h7FB56408A201;
			 12: q = 48'h7FA737096A90;
			 13: q = 48'h7F97CF0A3309;
			 14: q = 48'h7F872C0AFB68;
			 15: q = 48'h7F754E0BC3AC;
			 16: q = 48'h7F62370C8BD3;
			 17: q = 48'h7F4DE40D53DC;
			 18: q = 48'h7F38580E1BC3;
			 19: q = 48'h7F21920EE387;
			 20: q = 48'h7F09920FAB27;
			 21: q = 48'h7EF0581072A0;
			 22: q = 48'h7ED5E61139F1;
			 23: q = 48'h7EBA3A120117;
			 24: q = 48'h7E9D5612C810;
			 25: q = 48'h7E7F39138EDC;
			 26: q = 48'h7E5FE5145577;
			 27: q = 48'h7E3F58151BE0;
			 28: q = 48'h7E1D9415E214;
			 29: q = 48'h7DFA9916A813;
			 30: q = 48'h7DD667176DDA;
			 31: q = 48'h7DB0FE183367;
			 32: q = 48'h7D8A5F18F8B8;
			 33: q = 48'h7D628B19BDCC;
			 34: q = 48'h7D39811A82A0;
			 35: q = 48'h7D0F421B4733;
			 36: q = 48'h7CE3CF1C0B82;
			 37: q = 48'h7CB7271CCF8D;
			 38: q = 48'h7C894C1D9350;
			 39: q = 48'h7C5A3D1E56CA;
			 40: q = 48'h7C29FC1F19F9;
			 41: q = 48'h7BF8881FDCDC;
			 42: q = 48'h7BC5E3209F70;
			 43: q = 48'h7B920C2161B4;
			 44: q = 48'h7B5D042223A5;
			 45: q = 48'h7B26CB22E542;
			 46: q = 48'h7AEF6323A688;
			 47: q = 48'h7AB6CC246777;
			 48: q = 48'h7A7D0525280C;
			 49: q = 48'h7A421125E846;
			 50: q = 48'h7A05EF26A822;
			 51: q = 48'h79C89F27679E;
			 52: q = 48'h798A242826B9;
			 53: q = 48'h794A7C28E571;
			 54: q = 48'h7909A929A3C5;
			 55: q = 48'h78C7AC2A61B1;
			 56: q = 48'h7884842B1F35;
			 57: q = 48'h7840332BDC4E;
			 58: q = 48'h77FABA2C98FC;
			 59: q = 48'h77B4182D553B;
			 60: q = 48'h776C4F2E110A;
			 61: q = 48'h77235F2ECC68;
			 62: q = 48'h76D94A2F8752;
			 63: q = 48'h768E0F3041C7;
			 64: q = 48'h7641AF30FBC5;
			 65: q = 48'h75F42C31B54A;
			 66: q = 48'h75A586326E55;
			 67: q = 48'h7555BD3326E3;
			 68: q = 48'h7504D333DEF3;
			 69: q = 48'h74B2C9349682;
			 70: q = 48'h745F9E354D90;
			 71: q = 48'h740B5436041B;
			 72: q = 48'h73B5EC36BA20;
			 73: q = 48'h735F66376F9E;
			 74: q = 48'h7307C4382494;
			 75: q = 48'h72AF0638D8FF;
			 76: q = 48'h72552D398CDD;
			 77: q = 48'h71FA393A402E;
			 78: q = 48'h719E2D3AF2EF;
			 79: q = 48'h7141083BA51E;
			 80: q = 48'h70E2CC3C56BA;
			 81: q = 48'h7083793D07C2;
			 82: q = 48'h7023113DB833;
			 83: q = 48'h6FC1943E680B;
			 84: q = 48'h6F5F033F174A;
			 85: q = 48'h6EFB5F3FC5ED;
			 86: q = 48'h6E96AA4073F2;
			 87: q = 48'h6E30E3412159;
			 88: q = 48'h6DCA0D41CE1E;
			 89: q = 48'h6D6228427A42;
			 90: q = 48'h6CF9354325C1;
			 91: q = 48'h6C8F3543D09B;
			 92: q = 48'h6C2429447ACD;
			 93: q = 48'h6BB813452457;
			 94: q = 48'h6B4AF245CD36;
			 95: q = 48'h6ADCC9467568;
			 96: q = 48'h6A6D99471CED;
			 97: q = 48'h69FD6147C3C2;
			 98: q = 48'h698C244869E6;
			 99: q = 48'h6919E3490F58;
			100: q = 48'h68A69F49B415;
			101: q = 48'h6832584A581D;
			102: q = 48'h67BD104AFB6D;
			103: q = 48'h6746C84B9E04;
			104: q = 48'h66CF814C3FE0;
			105: q = 48'h66573D4CE100;
			106: q = 48'h65DDFC4D8163;
			107: q = 48'h6563C04E2106;
			108: q = 48'h64E8894EBFE9;
			109: q = 48'h646C5A4F5E09;
			110: q = 48'h63EF334FFB65;
			111: q = 48'h6371155097FC;
			112: q = 48'h62F2025133CD;
			113: q = 48'h6271FA51CED4;
			114: q = 48'h61F100526912;
			115: q = 48'h616F14530285;
			116: q = 48'h60EC38539B2B;
			117: q = 48'h60686D543302;
			118: q = 48'h5FE3B454CA0A;
			119: q = 48'h5F5E0E556041;
			120: q = 48'h5ED77D55F5A5;
			121: q = 48'h5E5001568A35;
			122: q = 48'h5DC79D571DEF;
			123: q = 48'h5D3E5257B0D2;
			124: q = 48'h5CB4215842DD;
			125: q = 48'h5C290B58D40F;
			126: q = 48'h5B9D11596465;
			127: q = 48'h5B103659F3DE;
			128: q = 48'h5A827A5A827A;
			129: q = 48'h59F3DE5B1036;
			130: q = 48'h5964655B9D11;
			131: q = 48'h58D40F5C290B;
			132: q = 48'h5842DD5CB421;
			133: q = 48'h57B0D25D3E52;
			134: q = 48'h571DEF5DC79D;
			135: q = 48'h568A355E5001;
			136: q = 48'h55F5A55ED77D;
			137: q = 48'h5560415F5E0E;
			138: q = 48'h54CA0A5FE3B4;
			139: q = 48'h54330260686D;
			140: q = 48'h539B2B60EC38;
			141: q = 48'h530285616F14;
			142: q = 48'h52691261F100;
			143: q = 48'h51CED46271FA;
			144: q = 48'h5133CD62F202;
			145: q = 48'h5097FC637115;
			146: q = 48'h4FFB6563EF33;
			147: q = 48'h4F5E09646C5A;
			148: q = 48'h4EBFE964E889;
			149: q = 48'h4E21066563C0;
			150: q = 48'h4D816365DDFC;
			151: q = 48'h4CE10066573D;
			152: q = 48'h4C3FE066CF81;
			153: q = 48'h4B9E046746C8;
			154: q = 48'h4AFB6D67BD10;
			155: q = 48'h4A581D683258;
			156: q = 48'h49B41568A69F;
			157: q = 48'h490F586919E3;
			158: q = 48'h4869E6698C24;
			159: q = 48'h47C3C269FD61;
			160: q = 48'h471CED6A6D99;
			161: q = 48'h4675686ADCC9;
			162: q = 48'h45CD366B4AF2;
			163: q = 48'h4524576BB813;
			164: q = 48'h447ACD6C2429;
			165: q = 48'h43D09B6C8F35;
			166: q = 48'h4325C16CF935;
			167: q = 48'h427A426D6228;
			168: q = 48'h41CE1E6DCA0D;
			169: q = 48'h4121596E30E3;
			170: q = 48'h4073F26E96AA;
			171: q = 48'h3FC5ED6EFB5F;
			172: q = 48'h3F174A6F5F03;
			173: q = 48'h3E680B6FC194;
			174: q = 48'h3DB833702311;
			175: q = 48'h3D07C2708379;
			176: q = 48'h3C56BA70E2CC;
			177: q = 48'h3BA51E714108;
			178: q = 48'h3AF2EF719E2D;
			179: q = 48'h3A402E71FA39;
			180: q = 48'h398CDD72552D;
			181: q = 48'h38D8FF72AF06;
			182: q = 48'h3824947307C4;
			183: q = 48'h376F9E735F66;
			184: q = 48'h36BA2073B5EC;
			185: q = 48'h36041B740B54;
			186: q = 48'h354D90745F9E;
			187: q = 48'h34968274B2C9;
			188: q = 48'h33DEF37504D3;
			189: q = 48'h3326E37555BD;
			190: q = 48'h326E5575A586;
			191: q = 48'h31B54A75F42C;
			192: q = 48'h30FBC57641AF;
			193: q = 48'h3041C7768E0F;
			194: q = 48'h2F875276D94A;
			195: q = 48'h2ECC6877235F;
			196: q = 48'h2E110A776C4F;
			197: q = 48'h2D553B77B418;
			198: q = 48'h2C98FC77FABA;
			199: q = 48'h2BDC4E784033;
			200: q = 48'h2B1F35788484;
			201: q = 48'h2A61B178C7AC;
			202: q = 48'h29A3C57909A9;
			203: q = 48'h28E571794A7C;
			204: q = 48'h2826B9798A24;
			205: q = 48'h27679E79C89F;
			206: q = 48'h26A8227A05EF;
			207: q = 48'h25E8467A4211;
			208: q = 48'h25280C7A7D05;
			209: q = 48'h2467777AB6CC;
			210: q = 48'h23A6887AEF63;
			211: q = 48'h22E5427B26CB;
			212: q = 48'h2223A57B5D04;
			213: q = 48'h2161B47B920C;
			214: q = 48'h209F707BC5E3;
			215: q = 48'h1FDCDC7BF888;
			216: q = 48'h1F19F97C29FC;
			217: q = 48'h1E56CA7C5A3D;
			218: q = 48'h1D93507C894C;
			219: q = 48'h1CCF8D7CB727;
			220: q = 48'h1C0B827CE3CF;
			221: q = 48'h1B47337D0F42;
			222: q = 48'h1A82A07D3981;
			223: q = 48'h19BDCC7D628B;
			224: q = 48'h18F8B87D8A5F;
			225: q = 48'h1833677DB0FE;
			226: q = 48'h176DDA7DD667;
			227: q = 48'h16A8137DFA99;
			228: q = 48'h15E2147E1D94;
			229: q = 48'h151BE07E3F58;
			230: q = 48'h1455777E5FE5;
			231: q = 48'h138EDC7E7F39;
			232: q = 48'h12C8107E9D56;
			233: q = 48'h1201177EBA3A;
			234: q = 48'h1139F17ED5E6;
			235: q = 48'h1072A07EF058;
			236: q = 48'h0FAB277F0992;
			237: q = 48'h0EE3877F2192;
			238: q = 48'h0E1BC37F3858;
			239: q = 48'h0D53DC7F4DE4;
			240: q = 48'h0C8BD37F6237;
			241: q = 48'h0BC3AC7F754E;
			242: q = 48'h0AFB687F872C;
			243: q = 48'h0A33097F97CF;
			244: q = 48'h096A907FA737;
			245: q = 48'h08A2017FB564;
			246: q = 48'h07D95C7FC256;
			247: q = 48'h0710A37FCE0C;
			248: q = 48'h0647D97FD888;
			249: q = 48'h057F007FE1C7;
			250: q = 48'h04B6197FE9CC;
			251: q = 48'h03ED277FF094;
			252: q = 48'h03242B7FF622;
			253: q = 48'h025B277FFA73;
			254: q = 48'h01921D7FFD88;
			255: q = 48'h00C9107FFF62;
			256: q = 48'h0000007FFFFF;
			257: q = 48'hFF36F07FFF62;
			258: q = 48'hFE6DE37FFD88;
			259: q = 48'hFDA4D97FFA73;
			260: q = 48'hFCDBD57FF622;
			261: q = 48'hFC12D97FF094;
			262: q = 48'hFB49E77FE9CC;
			263: q = 48'hFA81007FE1C7;
			264: q = 48'hF9B8277FD888;
			265: q = 48'hF8EF5D7FCE0C;
			266: q = 48'hF826A47FC256;
			267: q = 48'hF75DFF7FB564;
			268: q = 48'hF695707FA737;
			269: q = 48'hF5CCF77F97CF;
			270: q = 48'hF504987F872C;
			271: q = 48'hF43C547F754E;
			272: q = 48'hF3742D7F6237;
			273: q = 48'hF2AC247F4DE4;
			274: q = 48'hF1E43D7F3858;
			275: q = 48'hF11C797F2192;
			276: q = 48'hF054D97F0992;
			277: q = 48'hEF8D607EF058;
			278: q = 48'hEEC60F7ED5E6;
			279: q = 48'hEDFEE97EBA3A;
			280: q = 48'hED37F07E9D56;
			281: q = 48'hEC71247E7F39;
			282: q = 48'hEBAA897E5FE5;
			283: q = 48'hEAE4207E3F58;
			284: q = 48'hEA1DEC7E1D94;
			285: q = 48'hE957ED7DFA99;
			286: q = 48'hE892267DD667;
			287: q = 48'hE7CC997DB0FE;
			288: q = 48'hE707487D8A5F;
			289: q = 48'hE642347D628B;
			290: q = 48'hE57D607D3981;
			291: q = 48'hE4B8CD7D0F42;
			292: q = 48'hE3F47E7CE3CF;
			293: q = 48'hE330737CB727;
			294: q = 48'hE26CB07C894C;
			295: q = 48'hE1A9367C5A3D;
			296: q = 48'hE0E6077C29FC;
			297: q = 48'hE023247BF888;
			298: q = 48'hDF60907BC5E3;
			299: q = 48'hDE9E4C7B920C;
			300: q = 48'hDDDC5B7B5D04;
			301: q = 48'hDD1ABE7B26CB;
			302: q = 48'hDC59787AEF63;
			303: q = 48'hDB98897AB6CC;
			304: q = 48'hDAD7F47A7D05;
			305: q = 48'hDA17BA7A4211;
			306: q = 48'hD957DE7A05EF;
			307: q = 48'hD8986279C89F;
			308: q = 48'hD7D947798A24;
			309: q = 48'hD71A8F794A7C;
			310: q = 48'hD65C3B7909A9;
			311: q = 48'hD59E4F78C7AC;
			312: q = 48'hD4E0CB788484;
			313: q = 48'hD423B2784033;
			314: q = 48'hD3670477FABA;
			315: q = 48'hD2AAC577B418;
			316: q = 48'hD1EEF6776C4F;
			317: q = 48'hD1339877235F;
			318: q = 48'hD078AE76D94A;
			319: q = 48'hCFBE39768E0F;
			320: q = 48'hCF043B7641AF;
			321: q = 48'hCE4AB675F42C;
			322: q = 48'hCD91AB75A586;
			323: q = 48'hCCD91D7555BD;
			324: q = 48'hCC210D7504D3;
			325: q = 48'hCB697E74B2C9;
			326: q = 48'hCAB270745F9E;
			327: q = 48'hC9FBE5740B54;
			328: q = 48'hC945E073B5EC;
			329: q = 48'hC89062735F66;
			330: q = 48'hC7DB6C7307C4;
			331: q = 48'hC7270172AF06;
			332: q = 48'hC6732372552D;
			333: q = 48'hC5BFD271FA39;
			334: q = 48'hC50D11719E2D;
			335: q = 48'hC45AE2714108;
			336: q = 48'hC3A94670E2CC;
			337: q = 48'hC2F83E708379;
			338: q = 48'hC247CD702311;
			339: q = 48'hC197F56FC194;
			340: q = 48'hC0E8B66F5F03;
			341: q = 48'hC03A136EFB5F;
			342: q = 48'hBF8C0E6E96AA;
			343: q = 48'hBEDEA76E30E3;
			344: q = 48'hBE31E26DCA0D;
			345: q = 48'hBD85BE6D6228;
			346: q = 48'hBCDA3F6CF935;
			347: q = 48'hBC2F656C8F35;
			348: q = 48'hBB85336C2429;
			349: q = 48'hBADBA96BB813;
			350: q = 48'hBA32CA6B4AF2;
			351: q = 48'hB98A986ADCC9;
			352: q = 48'hB8E3136A6D99;
			353: q = 48'hB83C3E69FD61;
			354: q = 48'hB7961A698C24;
			355: q = 48'hB6F0A86919E3;
			356: q = 48'hB64BEB68A69F;
			357: q = 48'hB5A7E3683258;
			358: q = 48'hB5049367BD10;
			359: q = 48'hB461FC6746C8;
			360: q = 48'hB3C02066CF81;
			361: q = 48'hB31F0066573D;
			362: q = 48'hB27E9D65DDFC;
			363: q = 48'hB1DEFA6563C0;
			364: q = 48'hB1401764E889;
			365: q = 48'hB0A1F7646C5A;
			366: q = 48'hB0049B63EF33;
			367: q = 48'hAF6804637115;
			368: q = 48'hAECC3362F202;
			369: q = 48'hAE312C6271FA;
			370: q = 48'hAD96EE61F100;
			371: q = 48'hACFD7B616F14;
			372: q = 48'hAC64D560EC38;
			373: q = 48'hABCCFE60686D;
			374: q = 48'hAB35F65FE3B4;
			375: q = 48'hAA9FBF5F5E0E;
			376: q = 48'hAA0A5B5ED77D;
			377: q = 48'hA975CB5E5001;
			378: q = 48'hA8E2115DC79D;
			379: q = 48'hA84F2E5D3E52;
			380: q = 48'hA7BD235CB421;
			381: q = 48'hA72BF15C290B;
			382: q = 48'hA69B9B5B9D11;
			383: q = 48'hA60C225B1036;
			384: q = 48'hA57D865A827A;
			385: q = 48'hA4EFCA59F3DE;
			386: q = 48'hA462EF596465;
			387: q = 48'hA3D6F558D40F;
			388: q = 48'hA34BDF5842DD;
			389: q = 48'hA2C1AE57B0D2;
			390: q = 48'hA23863571DEF;
			391: q = 48'hA1AFFF568A35;
			392: q = 48'hA1288355F5A5;
			393: q = 48'hA0A1F2556041;
			394: q = 48'hA01C4C54CA0A;
			395: q = 48'h9F9793543302;
			396: q = 48'h9F13C8539B2B;
			397: q = 48'h9E90EC530285;
			398: q = 48'h9E0F00526912;
			399: q = 48'h9D8E0651CED4;
			400: q = 48'h9D0DFE5133CD;
			401: q = 48'h9C8EEB5097FC;
			402: q = 48'h9C10CD4FFB65;
			403: q = 48'h9B93A64F5E09;
			404: q = 48'h9B17774EBFE9;
			405: q = 48'h9A9C404E2106;
			406: q = 48'h9A22044D8163;
			407: q = 48'h99A8C34CE100;
			408: q = 48'h99307F4C3FE0;
			409: q = 48'h98B9384B9E04;
			410: q = 48'h9842F04AFB6D;
			411: q = 48'h97CDA84A581D;
			412: q = 48'h97596149B415;
			413: q = 48'h96E61D490F58;
			414: q = 48'h9673DC4869E6;
			415: q = 48'h96029F47C3C2;
			416: q = 48'h959267471CED;
			417: q = 48'h952337467568;
			418: q = 48'h94B50E45CD36;
			419: q = 48'h9447ED452457;
			420: q = 48'h93DBD7447ACD;
			421: q = 48'h9370CB43D09B;
			422: q = 48'h9306CB4325C1;
			423: q = 48'h929DD8427A42;
			424: q = 48'h9235F341CE1E;
			425: q = 48'h91CF1D412159;
			426: q = 48'h9169564073F2;
			427: q = 48'h9104A13FC5ED;
			428: q = 48'h90A0FD3F174A;
			429: q = 48'h903E6C3E680B;
			430: q = 48'h8FDCEF3DB833;
			431: q = 48'h8F7C873D07C2;
			432: q = 48'h8F1D343C56BA;
			433: q = 48'h8EBEF83BA51E;
			434: q = 48'h8E61D33AF2EF;
			435: q = 48'h8E05C73A402E;
			436: q = 48'h8DAAD3398CDD;
			437: q = 48'h8D50FA38D8FF;
			438: q = 48'h8CF83C382494;
			439: q = 48'h8CA09A376F9E;
			440: q = 48'h8C4A1436BA20;
			441: q = 48'h8BF4AC36041B;
			442: q = 48'h8BA062354D90;
			443: q = 48'h8B4D37349682;
			444: q = 48'h8AFB2D33DEF3;
			445: q = 48'h8AAA433326E3;
			446: q = 48'h8A5A7A326E55;
			447: q = 48'h8A0BD431B54A;
			448: q = 48'h89BE5130FBC5;
			449: q = 48'h8971F13041C7;
			450: q = 48'h8926B62F8752;
			451: q = 48'h88DCA12ECC68;
			452: q = 48'h8893B12E110A;
			453: q = 48'h884BE82D553B;
			454: q = 48'h8805462C98FC;
			455: q = 48'h87BFCD2BDC4E;
			456: q = 48'h877B7C2B1F35;
			457: q = 48'h8738542A61B1;
			458: q = 48'h86F65729A3C5;
			459: q = 48'h86B58428E571;
			460: q = 48'h8675DC2826B9;
			461: q = 48'h86376127679E;
			462: q = 48'h85FA1126A822;
			463: q = 48'h85BDEF25E846;
			464: q = 48'h8582FB25280C;
			465: q = 48'h854934246777;
			466: q = 48'h85109D23A688;
			467: q = 48'h84D93522E542;
			468: q = 48'h84A2FC2223A5;
			469: q = 48'h846DF42161B4;
			470: q = 48'h843A1D209F70;
			471: q = 48'h8407781FDCDC;
			472: q = 48'h83D6041F19F9;
			473: q = 48'h83A5C31E56CA;
			474: q = 48'h8376B41D9350;
			475: q = 48'h8348D91CCF8D;
			476: q = 48'h831C311C0B82;
			477: q = 48'h82F0BE1B4733;
			478: q = 48'h82C67F1A82A0;
			479: q = 48'h829D7519BDCC;
			480: q = 48'h8275A118F8B8;
			481: q = 48'h824F02183367;
			482: q = 48'h822999176DDA;
			483: q = 48'h82056716A813;
			484: q = 48'h81E26C15E214;
			485: q = 48'h81C0A8151BE0;
			486: q = 48'h81A01B145577;
			487: q = 48'h8180C7138EDC;
			488: q = 48'h8162AA12C810;
			489: q = 48'h8145C6120117;
			490: q = 48'h812A1A1139F1;
			491: q = 48'h810FA81072A0;
			492: q = 48'h80F66E0FAB27;
			493: q = 48'h80DE6E0EE387;
			494: q = 48'h80C7A80E1BC3;
			495: q = 48'h80B21C0D53DC;
			496: q = 48'h809DC90C8BD3;
			497: q = 48'h808AB20BC3AC;
			498: q = 48'h8078D40AFB68;
			499: q = 48'h8068310A3309;
			500: q = 48'h8058C9096A90;
			501: q = 48'h804A9C08A201;
			502: q = 48'h803DAA07D95C;
			503: q = 48'h8031F40710A3;
			504: q = 48'h8027780647D9;
			505: q = 48'h801E39057F00;
			506: q = 48'h80163404B619;
			507: q = 48'h800F6C03ED27;
			508: q = 48'h8009DE03242B;
			509: q = 48'h80058D025B27;
			510: q = 48'h80027801921D;
			511: q = 48'h80009E00C910;
		
		endcase
	end

endmodule

