module test(input btn, output led);
	assign led = btn;
endmodule