module sevenSegDisplay(
	/* TODO: Ports go here (refer to lab spec) */
);

	/* TODO: Instantiate six copies of sevenSegDigit, one for each digit (calculated below)*/

	// The following block will contain the logic of your combinational circuit
	always_comb begin
		/* TODO: Convert a 20-bit input number to six individual digits (4 bits each) */
	end

endmodule