module miniALU_top(input [9:0] switches, output [9:0] leds);
	
	assign leds = switches;
	

endmodule