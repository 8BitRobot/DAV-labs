module cube_top(
    input clk,
    output [15:0] M [0:3][0:3]
);
    reg [15:0] vertices [0:7][0:2] = '{'{0,0,0},'{0,0,1},'{0,1,0},'{0,1,1},'{1,0,0},'{1,0,1},'{1,1,0},'{1,1,1}};
    reg [15:0] indexed_face_set [0:11][0:2] = '{'{0,1,2},'{1,3,2},'{2,3,6},'{3,7,6},'{0,2,4},'{2,6,4},'{1,5,3},'{3,5,7},'{0,4,1},'{1,4,5},'{4,6,5},'{5,6,7}};
    
	 
	 
endmodule