module game_controller (
    input clk
);

endmodule
